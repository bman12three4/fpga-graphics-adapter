module ctxt_ctrl ();
endmodule
