module vga_ctrl (
		input vga_clk,
		
		output reg [9:0] posx,
		output reg [8:0] posy,
		
		output reg vsync,
		output reg hsync,
		
		output reg [9:0] h_pixel,
		output reg [9:0] line,
		
		input [3:0] r_in,
		input [3:0] g_in,
		input [3:0] b_in,
		
		output [3:0] r_out,
		output [3:0] g_out,
		output [3:0] b_out
	);
	

	end

	
endmodule
